----------------------------------------------------------------------------------
-- Projeto: processador simplificado
-- Modulo: registradores de dados - 1 entrada e 2 saidas.
-- Prof. Pedro L. Benko - FEI - 2011
-- 4 bits addrees; 8 bits data bus
-- regs.vhd
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--
entity regs is
	port (clock : in std_logic;
		  rst	: in std_logic;
		  RFwe	: in std_logic; -- enable escrita
		  RFr1e : in std_logic; -- enable leitura reg1
		  RFr2e	: in std_logic; -- enable leitura reg2
		  RFwa	: in std_logic_vector(3 downto 0);-- address escrita
		  RFr1a	: in std_logic_vector(3 downto 0);-- address leitura reg1
		  RFr2a	: in std_logic_vector(3 downto 0);-- address leitura reg2
		  RFw	: in std_logic_vector(7 downto 0);-- data escrita
		  RFr1	: out std_logic_vector(7 downto 0); -- data leitura reg1
		  RFr2	: out std_logic_vector(7 downto 0));-- data leitura reg2
end regs;
architecture behv of regs is
	type rf_type is array (0 to 15) of
	std_logic_vector(7 downto 0);
	signal tmp_rf: rf_type;
begin
----------------------------------------------------------------------------------
write: process(clock, rst, RFwa, RFwe, RFw)
begin
	if rst='0' then -- ativo em alto
		tmp_rf <= (tmp_rf'range => "00000000");
	else
		if (clock'event and clock = '1') then
			if RFwe='1' then
			tmp_rf(conv_integer(RFwa)) <= RFw;
			end if;
		end if;
	end if;
end process;
----------------------------------------------------------------------------------
read1: process(clock, rst, RFr1e, RFr1a)
begin
	if rst='0' then
	RFr1 <= "00000000";
	else
		if (clock'event and clock = '1') then
			if RFr1e='1' then
			RFr1 <= tmp_rf(conv_integer(RFr1a));
			end if;
		end if;
	end if;
end process;
----------------------------------------------------------------------------------
read2: process(clock, rst, RFr2e, RFr2a)
begin
	if rst='0' then
	RFr2<= "00000000";
	else
		if (clock'event and clock = '1') then
			if RFr2e='1' then
			RFr2 <= tmp_rf(conv_integer(RFr2a));
			end if;
		end if;
	end if;
end process;
end behv;
----------------------------------------------------------------------------------